class mimsg ;
  reg [31 :0] addr ;
  reg [31 :0] data ;
  reg rw ;
  
endclass 
